module control();



endmodule