module control();




endmodule