module onewire(in, out);
 
input in;
output out;


endmodule